package gap_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  typedef class gap_driver;
  typedef class gap_monitor;

  `include "gap_bfm_cb.svh"
  `include "gap_bfm.svh"

  `include "gap_base_cfg.svh"
  `include "gap_cfg.svh"

  `include "gap_driver.svh"
  `include "gap_monitor.svh"

  `include "gap_base_agent.svh"
  `include "gap_agent.svh"
endpackage : gap_pkg
